/*
 * Copyright (c) 2024 Tyler Hong
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_tyler_hong_onboarding (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    wire [7:0]  en_reg_out_7_0;
    wire [7:0]  en_reg_out_15_8;
    wire [7:0]  en_reg_pwm_7_0;
    wire [7:0]  en_reg_pwm_15_8;
    wire [7:0]  pwm_duty_cycle;
    wire [15:0] pwm_out;


    spi_peripheral spi_peripheral_instance (
        .clk              (clk),
        .rst_n            (rst_n),
        .ncs              (ui_in[2]),
        .sclk             (ui_in[0]),
        .copi             (ui_in[1]),
        .en_reg_out_7_0   (en_reg_out_7_0),
        .en_reg_out_15_8  (en_reg_out_15_8),
        .en_reg_pwm_7_0   (en_reg_pwm_7_0),
        .en_reg_pwm_15_8  (en_reg_pwm_15_8),
        .pwm_duty_cycle   (pwm_duty_cycle)
    );

    pwm_peripheral pwm_peripheral_instance (
        .clk              (clk),
        .rst_n            (rst_n),
        .en_reg_out_7_0   (en_reg_out_7_0),
        .en_reg_out_15_8  (en_reg_out_15_8),
        .en_reg_pwm_7_0   (en_reg_pwm_7_0),
        .en_reg_pwm_15_8  (en_reg_pwm_15_8),
        .pwm_duty_cycle   (pwm_duty_cycle),
        .out              (pwm_out)
    );

    assign uo_out  = pwm_out[7:0];
    assign uio_out = pwm_out[15:8];
    assign uio_oe  = 8'hFF;

    // List all unused inputs to prevent warnings.
    wire _unused = &{ena, ui_in[7:3], uio_in, 1'b0};

endmodule
